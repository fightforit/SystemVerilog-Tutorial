module mux_2to1 ();


endmodule : mux_2to1
