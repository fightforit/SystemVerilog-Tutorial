module mux_2to1 #(
    parameter int    BIT_WIDTH = 8,
    parameter string method    = "conti"
) (
    input  logic                 sel_i,
    input  logic [BIT_WIDTH-1:0] a_i,
    input  logic [BIT_WIDTH-1:0] b_i,
    output logic [BIT_WIDTH-1:0] y_o
);

  if (method == "conti") begin
    // Continuous assignment
    assign y_o = sel_i ? b_i : a_i;
  end else if (method == "proc1") begin
    // Procedural 1
    always_comb begin
      y_o = sel_i ? b_i : a_i;
    end
  end else if (method == "proc2") begin
    // Procedural 2
    always_comb begin
      if (sel_i) begin
        y_o = b_i;
      end else begin
        y_o = a_i;
      end
    end
  end

endmodule : mux_2to1
